package apb_slave_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "apb_slave_if.sv"
  `include "apb_slave_vif.sv"
  `include "apb_slave_seq_item.sv"
  `include "apb_slave_cfg.sv"
  `include "apb_slave_model.sv"
  `include "apb_slave_driver.sv"
  `include "apb_slave_monitor.sv"
  `include "apb_slave_agent.sv"
  `include "apb_slave_scoreboard.sv"
  `include "apb_slave_env.sv"
  `include "apb_slave_sequences.sv"

endpackage

