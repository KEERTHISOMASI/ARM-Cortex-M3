// ahb_master_sequencer.sv
`ifndef AHB_MASTER_SEQUENCER_SV
`define AHB_MASTER_SEQUENCER_SV 

typedef uvm_sequencer#(ahb_seq_item) ahb_master_sequencer;

`endif

