`ifndef AHB_SLAVE_SEQUENCER_SV
`define AHB_SLAVE_SEQUENCER_SV 

typedef uvm_sequencer#(ahb_seq_item) ahb_slave_sequencer;

`endif

