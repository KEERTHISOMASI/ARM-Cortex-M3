package sram_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "sram_if.sv"
  `include "sram_seq_item.sv"
  `include "sram_storage_c.sv"
  `include "sram_agent_config.sv"
  `include "sram_driver.sv"
  `include "sram_monitor.sv"
  `include "sram_agent.sv"

endpackage

