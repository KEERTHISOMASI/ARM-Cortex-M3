`ifndef APB_SLAVE_VIF_SV
`define APB_SLAVE_VIF_SV

typedef virtual apb_slave_if.slave_mp apb_slave_vif;

`endif

